(diagram:(two_terminal:[(((2,3),(2,1)),Battery(5.0)),(((1,1),(2,1)),Resistor(100.0)),(((1,3),(2,3)),Wire),(((1,0),(1,1)),Wire),(((1,0),(3,0)),Wire),(((3,0),(3,4)),Resistor(1000.0)),(((-1,4),(3,4)),Wire),(((-1,3),(-1,4)),Capacitor(0.0001)),(((-1,3),(-1,2)),Capacitor(0.0001)),(((-1,2),(0,2)),Wire),(((-2,4),(-2,2)),Inductor(0.08, None)),(((-1,3),(1,3)),Wire),(((-2,4),(-1,4)),Wire),(((-2,2),(-1,2)),Wire),(((2,3),(4,3)),Wire),(((2,1),(2,-1)),Wire),(((2,-1),(4,-1)),Wire),(((4,1),(4,3)),Resistor(1000.0)),(((5,0),(5,-1)),Wire),(((5,2),(5,3)),Resistor(10.0)),(((4,3),(5,3)),Wire),(((4,-1),(5,-1)),Wire)],three_terminal:[(((1,3),(0,2),(1,1)),NTransistor(100.0)),(((4,1),(3,0),(4,-1)),NTransistor(100.0)),(((5,2),(4,1),(5,0)),NTransistor(100.0))]),cfg:(max_nr_iters:200,nr_step_size:0.1,nr_tolerance:0.000000001,dx_soln_tolerance:0.001,mode:NewtonRaphson),dt:0.0001,sample_rate:6000)
