(diagram:(two_terminal:[(((1,4),(1,2)),Battery(5.0)),(((3,2),(3,4)),Inductor(1.0)),(((3,2),(5,2)),Capacitor(0.01)),(((5,2),(5,4)),Wire),(((1,4),(3,4)),Wire),(((1,2),(3,2)),Switch(false)),(((5,4),(3,4)),Capacitor(0.01)),(((5,4),(5,6)),Inductor(1.0)),(((3,6),(5,6)),Wire),(((3,4),(3,6)),Wire)],three_terminal:[]),cfg:(max_nr_iters:20,nr_step_size:0.1,nr_tolerance:0.001,dx_soln_tolerance:0.001,mode:Linear,adaptive_step_size:true,n_timesteps:2),dt:0.005,sample_rate:6000)
